
.subckt MAC8_24F 
+ w1_7 w1_6 w1_5 w1_4 w1_3 w1_2 w1_1 w1_0 							
+ w2_7 w2_6 w2_5 w2_4 w2_3 w2_2 w2_1 w2_0 
+ a7 a6 a5 a4 a3 a2 a1 a0  
+ b7 b6 b5 b4 b3 b2 b1 b0
+ z16 z15 z14 z13 z12 z11 z10 z9 z8 z7 z6 z5 z4 z3 z2 z1 z0


**********

.ends


*.subckt ***

***********

*.ends
