.subckt AN_lvt_2 A B out W=120n L=40n f=1
** TODO
.ends AN_lvt_2
