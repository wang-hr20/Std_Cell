.subckt OR_lvt_2 A B out W=120n L=40n f=1

.include ./NR_lvt_2.sp
.include ./Inv_lvt.sp

X_NR A B A_NR_B NR_lvt_2 f=f
X_Inv A_NR_B out Inv_lvt f=f
.ends OR_lvt_2
